----------------------------------------------------------------------------------
-- Company: THE Ohio State University
-- Engineer: Gage Farmer & Chloe Oh
-- 
-- Create Date:    14:48:33 03/28/2024 
-- Design Name: 	 System Controller
-- Module Name:    controller - Behavioral 
-- Project Name: 	 Project 3
-- Target Devices: Your mom
-- Tool versions:  14.7
-- Description:    It is a system controller mane
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity controller is
    Port ( CLK	: in STD_LOGIC;
			  M, N : in  STD_LOGIC_VECTOR (4 downto 1);
           ST : in  STD_LOGIC;
           DONE : out  STD_LOGIC;
			  R : out  STD_LOGIC_VECTOR (8 downto 1));
end controller;

entity shift_register is
		Port ( CLK	: in STD_LOGIC;
			  M, N : in  STD_LOGIC_VECTOR (4 downto 1);
           ST : in  STD_LOGIC;
           DONE : out  STD_LOGIC;
			  R : out  STD_LOGIC_VECTOR (8 downto 1));
end shift_register;

architecture Behavioral of controller is
	signal State: integer range 0 to 9;
	signal ACC: std_logic_vector(8 downto 0);		-- accumulator
	alias Z: std_logic is ACC(0);						-- Z is bit 0 of ACC
	
architecture Behavioural of shift_register is
	signal State:
	signal ACC:
	alias Z:
	
begin
		R <= ACC(7 downto 0);
		process (CLK)
		begin
			if CLK'event and CLK = '1' then			-- executes on rising edge
		
			case State is
			when 0 =>
				if ST = '1' then
					ACC(8 downto 4) <= "00000";		-- clear upper ACC
					ACC(3 downto 0) <= N;				-- load multiplier
					State <= 1;
				end if;
			when 1|3|5|7 =>								-- "add/shift" state
				if Z = '1' then							-- add multiplicand to ACC
					ACC(8 downto 4) <= ('0'&ACC(7 downto 4)) + M;
					State <= State + 1;
				else ACC <= '0'&ACC(8 downto 1);		-- shift accumulator right
					State <= State + 2;
				end if;
			when 2|4|6|8 =>								-- shift state
				ACC <= '0'&ACC(8 downto 1);			-- right shift
				State <= State + 1;
			when 9 =>										-- end of cycle
				State <= 0;
			end case;
			end if;
		end process;
		Done <= '1' when State = 9 else '0';


end Behavioral;

