library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Custom 9-bit Shift Register
entity custom_shift_reg is
  port (
    clk : in std_logic;
    S0, S1 : in std_logic;
    load, shift_right, shift_left : out std_logic;
    Q : buffer std_logic_vector(8 downto 0)
  );
end entity custom_shift_reg;

architecture behavioral of custom_shift_reg is
begin
  process (clk)
  begin
    if rising_edge(clk) then
      if S1 = '0' and S0 = '0' then
        load <= '1';
        shift_right <= '0';
        shift_left <= '0';
      elsif S1 = '0' and S0 = '1' then
        load <= '0';
        shift_right <= '1';
        shift_left <= '0';
      elsif S1 = '1' and S0 = '0' then
        load <= '0';
        shift_right <= '0';
        shift_left <= '1';
      elsif S1 = '1' and S0 = '1' then
        load <= '0';
        shift_right <= '0';
        shift_left <= '0';
      end if;
    end if;
  end process;
end architecture behavioral;

-- 4-bit Parallel Adder
entity parallel_adder is
  port (
    X, Y : in std_logic_vector(3 downto 0);
    C_in : in std_logic;
    sum : out std_logic_vector(3 downto 0);
    C_out : out std_logic
  );
end entity parallel_adder;

architecture behavioral of parallel_adder is
begin
  process (X, Y, C_in)
    variable temp_sum : std_logic_vector(4 downto 0);
  begin
    temp_sum := ('0' & X) + ('0' & Y) + C_in;
    sum <= temp_sum(3 downto 0);
    C_out <= temp_sum(4);
  end process;
end architecture behavioral;

-- System Controller
entity system_controller is
  port (
    clk, start : in std_logic;
    done : out std_logic
  );
end entity system_controller;

architecture behavioral of system_controller is
begin
  process (clk, start)
    variable state : integer := 0;
  begin
    if rising_edge(clk) then
      case state is
        when 0 =>
          if start = '1' then
            state := 1;
          end if;
        -- other states and transitions omitted for brevity
        when others =>
          state := 0;
      end case;
    end if;
    done <= '1' when state = 2 else '0';
  end process;
end architecture behavioral;

-- Multiplication Circuit
entity multiplier is
  port (
    clk, start : in std_logic;
    multiplicand, multiplier : in std_logic_vector(3 downto 0);
    result : out std_logic_vector(7 downto 0);
    done : out std_logic
  );
end entity multiplier;

architecture behavioral of multiplier is
  signal intermediate_result : std_logic_vector(7 downto 0) := (others => '0');
begin
  process (clk)
  begin
    if rising_edge(clk) then
      if start = '1' then
        intermediate_result <= (others => '0');
      elsif done = '0' then
        -- multiplication procedure
        -- logic to update intermediate_result based on multiplicand and multiplier
      end if;
    end if;
  end process;
  result <= intermediate_result;
end architecture behavioral;